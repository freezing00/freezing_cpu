LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY IR IS
PORT(
	D:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	CLK:IN STD_LOGIC;
	Q:OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END IR;
ARCHITECTURE A OF IR IS
BEGIN 
	PROCESS(CLK)
	BEGIN
		IF(CLK'EVENT AND CLK='1') THEN
			Q<=D;
		END IF;
	END PROCESS;
END A;
