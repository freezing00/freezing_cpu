LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY CONVERT IS
PORT(
     IRCODE:IN STD_LOGIC_VECTOR(15 DOWNTO 0);
	 OP:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
     I11,I10,I9,I8:OUT STD_LOGIC;
     A:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
	 );
END CONVERT;
ARCHITECTURE A OF CONVERT IS
BEGIN
   OP<=IRCODE(15 DOWNTO 12);
   I11<=IRCODE(11);
   I10<=IRCODE(10);
   I9<=IRCODE(9);
   I8<=IRCODE(8);
   A<=IRCODE(7 DOWNTO 0);
END A;
