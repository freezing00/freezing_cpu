LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY MUX4 IS
PORT(
	A,B:IN STD_LOGIC;
	X0,X1,X2,X3:IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	W:OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
);
END MUX4;
ARCHITECTURE A OF MUX4 IS
BEGIN
	PROCESS
	BEGIN
		IF(A='0'AND B='0')THEN
			W<=X0;
		ELSIF(A='0'AND B='1')THEN
			W<=X1;
		ELSIF(A='1'AND B='0')THEN
			W<=X2;
		ELSE
			W<=X3;
		END IF;
	END PROCESS;
END A;

