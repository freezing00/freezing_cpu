LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY MCOMMAND IS
PORT(
     T2,T3,T4:IN STD_LOGIC; 
     D:IN STD_LOGIC_VECTOR(20 DOWNTO 0);
     LOAD,LDPC,LDAR,LDIR,LDRI,LDPSW,RS_B,S2,S1,S0:OUT STD_LOGIC;
     ALU_B,SW_B,LED_B,RD_D,CS_D,RAM_B,CS_I,ADDR_B,P1,P2,p3:OUT STD_LOGIC        
    );
END  MCOMMAND;
ARCHITECTURE A OF MCOMMAND IS
SIGNAL DATAOUT:STD_LOGIC_VECTOR(20 DOWNTO 0);
BEGIN 
PROCESS(T2,T3,T4,DATAOUT)
    BEGIN
        IF(T2'EVENT AND T2='1') THEN
             DATAOUT(20 DOWNTO 0)<=D(20 DOWNTO 0);
        END IF;
		LOAD<=DATAOUT(20);
		LDPC<=DATAOUT(19) AND T4;
		LDAR<=DATAOUT(18) AND T3;
		LDIR<=DATAOUT(17) AND T3;
		LDRI<=DATAOUT(16) AND T4;
		LDPSW<=DATAOUT(15) AND T3;
		RS_B<=DATAOUT(14);
		S2<=DATAOUT(13);
		S1<=DATAOUT(12);
		S0<=DATAOUT(11);
		ALU_B<=DATAOUT(10);
		SW_B<=DATAOUT(9);
		LED_B<=DATAOUT(8);
		RD_D<=DATAOUT(7);
		CS_D<=DATAOUT(6)AND T3;
		RAM_B<=DATAOUT(5);
		CS_I<=DATAOUT(4);
		ADDR_B<=DATAOUT(3);
		P1<=DATAOUT(2);
		P2<=DATAOUT(1);
		P3<=DATAOUT(0);
    END PROCESS;
END A;


